library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

entity InstructionMemory is
    Port ( I_clk : in  STD_LOGIC;
           I_addr : in  STD_LOGIC_VECTOR (15 downto 0);
           O_data : out  STD_LOGIC_VECTOR (31 downto 0));
end InstructionMemory;

architecture Behavioral of InstructionMemory is
	type store_t is array (0 to 255) of std_logic_vector(31 downto 0);
   signal InstructionMemory: store_t := (
		--0 => "00000000111001110000100000100000", -- add
		--1 => "00000000111001010001000000100010", -- subtract
		--2 => "00000000001000100001100000100100", -- and
		--3 => "00000000001000100010000000100101", -- or
		--4 => "00000000001000100010100000100110", --- xor
      --5 => "00000000001000100011000000100111", --- nor
		--6 => "00000000011000100011100000101010", --- slt
		--7 => "00000000110000100001000000101001", --- sltu
		--8 => "00000000000000010011100101000000", --- sll
		--9 => "00000000000000010011000101000010", --- srl
		--10 =>"00000000000001000010100101000011", --- sra
		--11 =>"00000000001000110010000000000100", --- sllv 
		--12 =>"00000000001001100001100000000110", --- srlv
		--13 =>"00000000111001010001000000000111", --- srav
		--14 =>"00000000110001010000100000100001", --- addu
		--15 =>"00000000010000010001100000100011", --- subu
		--16 => "10001100001000100000000000000100", -- lw  $2, 4($1)
		--17 => "10000000001000110000000000000101", -- lb  $3, 5($1)
		--18 => "10000100001001000000000000001000", -- lh  $4, 8($1)
		--19 => "10010000001001010000000000001100", -- lbu $5, 12($1)
		--20 => "10010100001001100000000000010000", -- lhu $6, 16($1)
		
		--0 => "10001100001000100000000000000100", -- lw  $2, 4($1)
		--1 => "10000000001000110000000000000111", -- lb  $3, 7($1)
		--2 => "10000100001001000000000000001000", -- lh  $4, 8($1)
		--3 => "10010000001001010000000000001100", -- lbu $5, 12($1)
		--4 => "10010100001001100000000000010000",  -- lhu $6, 16($1)
		
		--5 => "10101100001001110000000000010100", -- sw $7, 20($1)
		--6 => "10100100001010000000000000010110", -- sh $8, 22($1)
		--7 => "10100000001010010000000000011000", -- sb $9, 24($1)
		
		--0 => "00100000000000010000000000001010", -- addi $1, $0, 10
		--1 => "00100000001000100000000000010100", -- addiu $2, $1, 20
		--2 => "00101000010000110000000000110010", -- slti $3, $2, 50
		--3 => "00101100010001000000000000001010", -- sltiu $4, $2, 10
		--4 => "00110000010001010000000000001111", -- andi $5, $2, 15
		--5 => "00110100010001100000000000000101", -- ori $6, $2, 5
		--6 => "00111000010001110000000000011001", -- xori $7, $2, 25
		--7 => "00111100000000100001001000110100", -- lui $2, 0x1234
		
		 --0  => "00100000000000010000000000000101",  -- addi $1, $0, 5     → $1 = 5
		 --1  => "00000000000000000000000000000000",  -- nop
		 --2  => "00000000000000000000000000000000",  -- nop
		 --3  => "00000000000000000000000000000000",  -- nop
		 
		 --4  => "00100000001000100000000000000011",  -- addi $2, $1, 3     → $2 = 8
		 --5  => "00000000000000000000000000000000",  -- nop
		 --6  => "00000000000000000000000000000000",  -- nop
		 --7  => "00000000000000000000000000000000",  -- nop
		 
		 --8  => "00100000000001000000000001010001",  -- addi $4, $0, 81    → $4 = 0x51
		 --9  => "00000000000000000000000000000000",  -- nop
		 --10 => "00000000000000000000000000000000",  -- nop
		 --11 => "00000000000000000000000000000000",  -- nop
		 
		 --12 => "00100000000001010000000000011001",  -- addi $5, $0, 25    → $5 = 0x19
		 --13 => "00000000000000000000000000000000",  -- nop
		 --14 => "00000000000000000000000000000000",  -- nop
		 --15 => "00000000000000000000000000000000",  -- nop
		 
		 --16 => "00100000000001100000000000010100",  -- addi $6, $0, 20    → $6 = 0x14
		 --17 => "00000000000000000000000000000000",  -- nop
		 --18 => "00000000000000000000000000000000",  -- nop
		 --19 => "00000000000000000000000000000000",  -- nop
		 
		 --20 => "00100000000001110000000000011011",  -- addi $7, $0, 27    → $7 = 0x1B
		 --21 => "00000000000000000000000000000000",  -- nop
		 --22 => "00000000000000000000000000000000",  -- nop
		 --23 => "00000000000000000000000000000000",  -- nop
		 
		 --24 => "00001000000000000000000000011000",  -- j 24 (infinite loop)
		 
    -- ==========================================
    -- SETUP: Initialize registers
    -- ==========================================
	--0  => x"20010005", -- addi  $1, $0, 5      ; $1 = 5
  	--1  => x"20030007", -- addi  $3, $0, 7      ; $3 = 7

  	-- EX -> EX forwarding: producer at 2, consumer at 3 (no NOP)
  	--2  => x"00231020", -- add   $2, $1, $3     ; $2 = $1 + $3 = 12
  	--3  => x"00432020", -- add   $4, $2, $3     ; $4 = $2 + $3 = 19 (EX->EX forward)

  	-- Mix of EX/MEM and MEM/WB forwarding
  	--4  => x"00233020", -- add   $6, $1, $3     ; $6 = $1 + $3 = 12
  	--5  => x"00C22820", -- add   $5, $6, $2     ; $5 = $6 + $2 = 24

  	-- Overwrite and forward to both inputs
  	--6  => x"00211020", -- add   $2, $1, $1     ; $2 = $1 + $1 = 10
  	--7  => x"00422020", -- add   $4, $2, $2     ; $4 = $2 + $2 = 20

  	-- Store & Load: no store->load bypass in your design, so insert NOP between SW and LW
  	--8  => x"AC020000", -- sw    $2, 0($0)      ; store $2 (10) to memory[0]
  	--9  => x"00000000", -- nop                  ; ensure store commits
 	--10  => x"8C020000", -- lw    $2, 0($0)      ; load $2 <= memory[0]
 	--11  => x"00000000", -- nop                  ; ensure load data available (load-use)

 	--12 => x"00432820", -- add   $5, $2, $3      ; $5 = $2 + $3 = 10 + 7 = 17
 	--13 => x"00443020", -- add   $6, $2, $4      ; $6 = $2 + $4 = 10 + 20 = 30

 	-- Branch operand forwarding test (producer at 16, BEQ at 17 uses forwarded value)
 	--14 => x"20010004", -- addi  $1, $0, 4      ; $1 = 4
 	--15 => x"20030004", -- addi  $3, $0, 4      ; $3 = 4
 	--16 => x"00201020", -- add   $2, $1, $0     ; $2 = $1 (copy $1 -> $2)
 	--17 => x"10430001", -- beq   $2, $3, +1     ; if $2 == $3 branch to addr 19 (tests branch forwarding)
 	--18 => x"20070001", -- addi  $7, $0, 1      ; not-taken path -> $7 = 1
 	--19 => x"20070002", -- addi  $7, $0, 2      ; taken path -> $7 = 2 (should execute when branch taken)

 	-- JR forwarding test: target produced by previous instruction (uses forwardedA)
 	--20 => x"20020017", -- addi  $2, $0, 23     ; FIXED: set $2 = 23 (instruction index)
 	--21 => x"00400008", -- jr    $2             ; jump to addr 23
 	--22 => x"20030001", -- addi  $3, $0, 1      ; skipped if JR worked
 	--23 => x"20030002", -- addi  $3, $0, 2      ; target: $3 = 2
	--24 => x"08000018", -- j     24             ; HALT: jump to self (infinite loop)
	0  => x"20010004", -- addi  $1, $0, 4      ; $1 = 4
	1  => x"20020004", -- addi  $2, $0, 4      ; $2 = 4
	2  => x"10220001", -- beq   $1, $2, +1     ; TAKEN (should predict correctly after first run)
	3  => x"20030001", -- addi  $3, $0, 1      ; SKIPPED
	4  => x"20030002", -- addi  $3, $0, 2      ; EXECUTED
	5  => x"08000000", -- j     0              ; Loop back to test prediction
	others => (others => '0')
		);
begin

	--process (I_clk)
	--begin
		--if rising_edge(I_clk) then
			--O_data <= InstructionMemory(to_integer(unsigned(I_addr(5 downto 0))));
		--end if;
	--end process;
	O_data <= InstructionMemory(to_integer(unsigned(I_addr(7 downto 0))));
end Behavioral;